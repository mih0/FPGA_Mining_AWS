/*
 * Copyright (c) 2017 Sprocket
 *
 * This is free software: you can redistribute it and/or modify
 * it under the terms of the GNU Affero General Public License with
 * additional permissions to the one published by the Free Software
 * Foundation, either version 3 of the License, or (at your option)
 * any later version. For more information see LICENSE.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Affero General Public License for more details.
 *
 * You should have received a copy of the GNU Affero General Public License
 * along with this program. If not, see <http://www.gnu.org/licenses/>.
 */

module fugue512 (
	input clk,
	input [511:0] data,
	output [511:0] hash
);
	
	reg [1151:0] S0, S1, S2, S3, S4, S5, S6, S7, S8;
	reg [1151:0] S9,S10,S11,S12,S13,S14,S15,S16,S17,S18;
	
	reg [511:0] H;
	
	assign hash = H;

	reg [511:0] x0, x0_1, x0_2, x0_3, x0_4, x0_5;
	reg [479:0] x1, x1_1, x1_2, x1_3, x1_4, x1_5;
	reg [447:0] x2, x2_1, x2_2, x2_3, x2_4, x2_5;
	reg [415:0] x3, x3_1, x3_2, x3_3, x3_4, x3_5;
	reg [383:0] x4, x4_1, x4_2, x4_3, x4_4, x4_5;
	reg [351:0] x5, x5_1, x5_2, x5_3, x5_4, x5_5;
	reg [319:0] x6, x6_1, x6_2, x6_3, x6_4, x6_5;
	reg [287:0] x7, x7_1, x7_2, x7_3, x7_4, x7_5;
	reg [255:0] x8, x8_1, x8_2, x8_3, x8_4, x8_5;
	reg [223:0] x9, x9_1, x9_2, x9_3, x9_4, x9_5;
	reg [191:0] x10, x10_1, x10_2, x10_3, x10_4, x10_5;
	reg [159:0] x11, x11_1, x11_2, x11_3, x11_4, x11_5;
	reg [127:0] x12, x12_1, x12_2, x12_3, x12_4, x12_5;
	reg [ 95:0] x13, x13_1, x13_2, x13_3, x13_4, x13_5;
	reg [ 63:0] x14, x14_1, x14_2, x14_3, x14_4, x14_5;
	reg [ 31:0] x15, x15_1, x15_2, x15_3, x15_4, x15_5;

	wire [1151:0] S1_d, S2_d, S3_d, S4_d, S5_d, S6_d, S7_d;
	wire [1151:0] S8_d, S9_d, S10_d, S11_d, S12_d, S13_d, S14_d, S15_d, S16_d, S17_d, S18_d;

	wire [1151:0] C0,C1,C2,C3,C4,C5,C6,C7;
	wire [1151:0] C8,C9,C10,C11,C12,C13,C14,C15;
	wire [1151:0] C16,C17,C18,C19,C20,C21,C22,C23;
	wire [1151:0] C24,C25,C26,C27,C28,C29,C30,C31,C32;	

	wire [1151:0] D0,D1,D2,D3,D4,D5,D6,D7;
	wire [1151:0] D8,D9,D10,D11,D12;
	
	round r0  (clk, x0[511:480], S0,  S1_d);
	round r1  (clk, x1[479:448], S1,  S2_d);
	round r2  (clk, x2[447:416], S2,  S3_d);
	round r3  (clk, x3[415:384], S3,  S4_d);
	round r4  (clk, x4[383:352], S4,  S5_d);
	round r5  (clk, x5[351:320], S5,  S6_d);
	round r6  (clk, x6[319:288], S6,  S7_d);
	round r7  (clk, x7[287:256], S7,  S8_d);
	round r8  (clk, x8[255:224], S8,  S9_d);
	round r9  (clk, x9[223:192], S9,  S10_d);
	round r10 (clk, x10[191:160], S10, S11_d);
	round r11 (clk, x11[159:128], S11, S12_d);
	round r12 (clk, x12[127: 96], S12, S13_d);
	round r13 (clk, x13[ 95: 64], S13, S14_d);
	round r14 (clk, x14[ 63: 32], S14, S15_d);
	round r15 (clk, x15[ 31:  0], S15, S16_d);
	round r16 (clk, 32'h00000000,  S16, S17_d);
	round r17 (clk, 32'h00000200,  S17, S18_d);
	
	close_1 c0 (clk, S18, C0);
	close_1 c1 (clk, C0, C1);
	close_1 c2 (clk, C1, C2);
	close_1 c3 (clk, C2, C3);
	close_1 c4 (clk, C3, C4);
	close_1 c5 (clk, C4, C5);
	close_1 c6 (clk, C5, C6);
	close_1 c7 (clk, C6, C7);
	close_1 c8 (clk, C7, C8);
	close_1 c9 (clk, C8, C9);
	close_1 c10 (clk, C9, C10);
	close_1 c11 (clk, C10, C11);
	close_1 c12 (clk, C11, C12);
	close_1 c13 (clk, C12, C13);
	close_1 c14 (clk, C13, C14);
	close_1 c15 (clk, C14, C15);
	close_1 c16 (clk, C15, C16);
	close_1 c17 (clk, C16, C17);
	close_1 c18 (clk, C17, C18);
	close_1 c19 (clk, C18, C19);
	close_1 c20 (clk, C19, C20);
	close_1 c21 (clk, C20, C21);
	close_1 c22 (clk, C21, C22);
	close_1 c23 (clk, C22, C23);
	close_1 c24 (clk, C23, C24);
	close_1 c25 (clk, C24, C25);
	close_1 c26 (clk, C25, C26);
	close_1 c27 (clk, C26, C27);
	close_1 c28 (clk, C27, C28);
	close_1 c29 (clk, C28, C29);
	close_1 c30 (clk, C29, C30);
	close_1 c31 (clk, C30, C31);

	close_2 d0 (clk, C31, D0);
	close_2 d1 (clk, D0, D1);
	close_2 d2 (clk, D1, D2);
	close_2 d3 (clk, D2, D3);
	close_2 d4 (clk, D3, D4);
	close_2 d5 (clk, D4, D5);
	close_2 d6 (clk, D5, D6);
	close_2 d7 (clk, D6, D7);
	close_2 d8 (clk, D7, D8);
	close_2 d9 (clk, D8, D9);
	close_2 d10 (clk, D9, D10);
	close_2 d11 (clk, D10, D11);
	close_2 d12 (clk, D11, D12);
	
	always @ (posedge clk) begin

			S0[1151:640] = 512'he13e3567da6ed11d951fddd625ea78e7437f203fcae65838ddb21398aac6e2c94a92efd106e8020bb6eecc54d915f117ac9ab027c5d3e4dbe616af758807a57e;
			S0[639:0] = 640'd0;
			
			S1 = { S1_d[767:0], S1_d[1151:768] };
			S2 = { S2_d[767:0], S2_d[1151:768] };
			S3 = { S3_d[767:0], S3_d[1151:768] };
			S4 = { S4_d[767:0], S4_d[1151:768] };
			S5 = { S5_d[767:0], S5_d[1151:768] };
			S6 = { S6_d[767:0], S6_d[1151:768] };
			S7 = { S7_d[767:0], S7_d[1151:768] };
			S8 = { S8_d[767:0], S8_d[1151:768] };
			S9 = { S9_d[767:0], S9_d[1151:768] };
			S10 = { S10_d[767:0], S10_d[1151:768] };
			S11 = { S11_d[767:0], S11_d[1151:768] };
			S12 = { S12_d[767:0], S12_d[1151:768] };
			S13 = { S13_d[767:0], S13_d[1151:768] };
			S14 = { S14_d[767:0], S14_d[1151:768] };
			S15 = { S15_d[767:0], S15_d[1151:768] };
			S16 = { S16_d[767:0], S16_d[1151:768] };
			S17 = { S17_d[767:0], S17_d[1151:768] };
			S18 = { S18_d[767:0], S18_d[1151:768] };
			
//			$display("S15: %x", S15[1151:640]);
//			$display("S18: %x", S18[1151:640]);
//			$display("C31: %x", C31[1151:640]);
//			$display("C31: %x", C31);
//			$display("D12: %x", D12[1151:640]);

			H = { D12[ 32 +: 32],
					D12[ 64 +: 32],
					D12[ 96 +: 32],
					D12[128 +: 32] ^ D12[0 +: 32],
					D12[288 +: 32] ^ D12[0 +: 32],
					D12[320 +: 32],
					D12[352 +: 32],
					D12[384 +: 32],
					D12[576 +: 32] ^ D12[0 +: 32],
					D12[608 +: 32],
					D12[640 +: 32],
					D12[672 +: 32],
					D12[864 +: 32] ^ D12[0 +: 32],
					D12[896 +: 32],
					D12[928 +: 32],
					D12[960 +: 32] };

		x15 = x15_5;
		x15_5 = x15_4;
		x15_4 = x15_3;
		x15_3 = x15_2;
		x15_2 = x15_1;
		x15_1 = x14[31:0];
		x14 = x14_5;
		x14_5 = x14_4;
		x14_4 = x14_3;
		x14_3 = x14_2;
		x14_2 = x14_1;
		x14_1 = x13[63:0];
		x13 = x13_5;
		x13_5 = x13_4;
		x13_4 = x13_3;
		x13_3 = x13_2;
		x13_2 = x13_1;
		x13_1 = x12[95:0];
		x12 = x12_5;
		x12_5 = x12_4;
		x12_4 = x12_3;
		x12_3 = x12_2;
		x12_2 = x12_1;
		x12_1 = x11[127:0];
		x11 = x11_5;
		x11_5 = x11_4;
		x11_4 = x11_3;
		x11_3 = x11_2;
		x11_2 = x11_1;
		x11_1 = x10[159:0];
		x10 = x10_5;
		x10_5 = x10_4;
		x10_4 = x10_3;
		x10_3 = x10_2;
		x10_2 = x10_1;
		x10_1 = x9[191:0];
		x9 = x9_5;
		x9_5 = x9_4;
		x9_4 = x9_3;
		x9_3 = x9_2;
		x9_2 = x9_1;
		x9_1 = x8[223:0];
		x8 = x8_5;
		x8_5 = x8_4;
		x8_4 = x8_3;
		x8_3 = x8_2;
		x8_2 = x8_1;
		x8_1 = x7[255:0];
		x7 = x7_5;
		x7_5 = x7_4;
		x7_4 = x7_3;
		x7_3 = x7_2;
		x7_2 = x7_1;
		x7_1 = x6[287:0];
		x6 = x6_5;
		x6_5 = x6_4;
		x6_4 = x6_3;
		x6_3 = x6_2;
		x6_2 = x6_1;
		x6_1 = x5[319:0];
		x5 = x5_5;
		x5_5 = x5_4;
		x5_4 = x5_3;
		x5_3 = x5_2;
		x5_2 = x5_1;
		x5_1 = x4[351:0];
		x4 = x4_5;
		x4_5 = x4_4;
		x4_4 = x4_3;
		x4_3 = x4_2;
		x4_2 = x4_1;
		x4_1 = x3[383:0];
		x3 = x3_5;
		x3_5 = x3_4;
		x3_4 = x3_3;
		x3_3 = x3_2;
		x3_2 = x3_1;
		x3_1 = x2[415:0];
		x2 = x2_5;
		x2_5 = x2_4;
		x2_4 = x2_3;
		x2_3 = x2_2;
		x2_2 = x2_1;
		x2_1 = x1[447:0];
		x1 = x1_5;
		x1_5 = x1_4;
		x1_4 = x1_3;
		x1_3 = x1_2;
		x1_2 = x1_1;
		x1_1 = x0[479:0];
		x0 = x0_5;
		x0_5 = x0_4;
		x0_4 = x0_3;
		x0_3 = x0_2;
		x0_2 = x0_1;
		x0_1 = data;
		
//		$display("S14:  %x", S14[1151:640]);
//		$display("x15:  %x", x15[ 31:  0]);
//		$display("S15x: %x", S15_d);
//		$display("S15:  %x", S15[1151:640]);
//		$display("S16x: %x", S16_d);

	end

endmodule

module round (
	input clk,
	input [31:0] q,
	input [1151:0] S,
	output [1151:0] O
);

	wire [127:0] S1, S2, S3, S4;

	reg [1151:0] S0_d, S1_d, S2_d, S3_d, S4_d;
	reg [1151:0] S0_q, S1_q, S2_q, S3_q, S4_q;
	
	smix smix0(S0_q[1152-((36-33)*32) +: 32], S0_q[1152-((36-34)*32) +: 32], S0_q[1152-((36-35)*32) +: 32], S0_q[1152-((36- 0)*32) +: 32], S1);
	smix smix1(S1_q[1152-((36-30)*32) +: 32], S1_q[1152-((36-31)*32) +: 32], S1_q[1152-((36-32)*32) +: 32], S1_q[1152-((36-33)*32) +: 32], S2);
	smix smix2(S2_q[1152-((36-27)*32) +: 32], S2_q[1152-((36-28)*32) +: 32], S2_q[1152-((36-29)*32) +: 32], S2_q[1152-((36-30)*32) +: 32], S3);
	smix smix3(S3_q[1152-((36-24)*32) +: 32], S3_q[1152-((36-25)*32) +: 32], S3_q[1152-((36-26)*32) +: 32], S3_q[1152-((36-27)*32) +: 32], S4);
	
	assign O = S4_q;
	
	always @ (*) begin
	
		S0_d = S;

		// TIX4
		S0_d[1152-((36-22)*32) +: 32] = S0_d[1152-((36-22)*32) +: 32] ^ S0_d[1152-((36- 0)*32) +: 32];
		S0_d[1152-((36- 0)*32) +: 32] = q;
		S0_d[1152-((36- 8)*32) +: 32] = S0_d[1152-((36- 8)*32) +: 32] ^ S0_d[1152-((36- 0)*32) +: 32];
		S0_d[1152-((36- 1)*32) +: 32] = S0_d[1152-((36- 1)*32) +: 32] ^ S0_d[1152-((36-24)*32) +: 32];
		S0_d[1152-((36- 4)*32) +: 32] = S0_d[1152-((36- 4)*32) +: 32] ^ S0_d[1152-((36-27)*32) +: 32];
		S0_d[1152-((36- 7)*32) +: 32] = S0_d[1152-((36- 7)*32) +: 32] ^ S0_d[1152-((36-30)*32) +: 32];

		// CMIX36 - 1
		S0_d[1152-((36-33)*32) +: 32] = S0_d[1152-((36-33)*32) +: 32] ^ S0_d[1152-((36- 1)*32) +: 32];
		S0_d[1152-((36-34)*32) +: 32] = S0_d[1152-((36-34)*32) +: 32] ^ S0_d[1152-((36- 2)*32) +: 32];
		S0_d[1152-((36-35)*32) +: 32] = S0_d[1152-((36-35)*32) +: 32] ^ S0_d[1152-((36- 3)*32) +: 32];
		S0_d[1152-((36-15)*32) +: 32] = S0_d[1152-((36-15)*32) +: 32] ^ S0_d[1152-((36- 1)*32) +: 32];
		S0_d[1152-((36-16)*32) +: 32] = S0_d[1152-((36-16)*32) +: 32] ^ S0_d[1152-((36- 2)*32) +: 32];
		S0_d[1152-((36-17)*32) +: 32] = S0_d[1152-((36-17)*32) +: 32] ^ S0_d[1152-((36- 3)*32) +: 32];
		
		S1_d = S0_q;
		S1_d[1087:1056] = S1[127:96];
		S1_d[1119:1088] = S1[95:64];
		S1_d[1151:1120] = S1[63:32];
		S1_d[31:0] = S1[31:0];

		// CMIX36 - 2
		S1_d[1152-((36-30)*32) +: 32] = S1_d[1152-((36-30)*32) +: 32] ^ S1_d[1152-((36-34)*32) +: 32];
		S1_d[1152-((36-31)*32) +: 32] = S1_d[1152-((36-31)*32) +: 32] ^ S1_d[1152-((36-35)*32) +: 32];
		S1_d[1152-((36-32)*32) +: 32] = S1_d[1152-((36-32)*32) +: 32] ^ S1_d[1152-((36- 0)*32) +: 32];
		S1_d[1152-((36-12)*32) +: 32] = S1_d[1152-((36-12)*32) +: 32] ^ S1_d[1152-((36-34)*32) +: 32];
		S1_d[1152-((36-13)*32) +: 32] = S1_d[1152-((36-13)*32) +: 32] ^ S1_d[1152-((36-35)*32) +: 32];
		S1_d[1152-((36-14)*32) +: 32] = S1_d[1152-((36-14)*32) +: 32] ^ S1_d[1152-((36- 0)*32) +: 32];

		S2_d = S1_q;
		S2_d[ 991:960] = S2[127:96];
		S2_d[1023:992] = S2[95:64];
		S2_d[1055:1024] = S2[63:32];
		S2_d[1087:1056] = S2[31:0];

		// CMIX36 - 3
		S2_d[1152-((36-27)*32) +: 32] = S2_d[1152-((36-27)*32) +: 32] ^ S2_d[1152-((36-31)*32) +: 32];
		S2_d[1152-((36-28)*32) +: 32] = S2_d[1152-((36-28)*32) +: 32] ^ S2_d[1152-((36-32)*32) +: 32];
		S2_d[1152-((36-29)*32) +: 32] = S2_d[1152-((36-29)*32) +: 32] ^ S2_d[1152-((36-33)*32) +: 32];
		S2_d[1152-((36- 9)*32) +: 32] = S2_d[1152-((36- 9)*32) +: 32] ^ S2_d[1152-((36-31)*32) +: 32];
		S2_d[1152-((36-10)*32) +: 32] = S2_d[1152-((36-10)*32) +: 32] ^ S2_d[1152-((36-32)*32) +: 32];
		S2_d[1152-((36-11)*32) +: 32] = S2_d[1152-((36-11)*32) +: 32] ^ S2_d[1152-((36-33)*32) +: 32];

		S3_d = S2_q;
		S3_d[895:864] = S3[127:96];
		S3_d[927:896] = S3[95:64];
		S3_d[959:928] = S3[63:32];
		S3_d[991:960] = S3[31:0];
		
		// CMIX36 - 4
		S3_d[1152-((36-24)*32) +: 32] = S3_d[1152-((36-24)*32) +: 32] ^ S3_d[1152-((36-28)*32) +: 32];
		S3_d[1152-((36-25)*32) +: 32] = S3_d[1152-((36-25)*32) +: 32] ^ S3_d[1152-((36-29)*32) +: 32];
		S3_d[1152-((36-26)*32) +: 32] = S3_d[1152-((36-26)*32) +: 32] ^ S3_d[1152-((36-30)*32) +: 32];
		S3_d[1152-((36- 6)*32) +: 32] = S3_d[1152-((36- 6)*32) +: 32] ^ S3_d[1152-((36-28)*32) +: 32];
		S3_d[1152-((36- 7)*32) +: 32] = S3_d[1152-((36- 7)*32) +: 32] ^ S3_d[1152-((36-29)*32) +: 32];
		S3_d[1152-((36- 8)*32) +: 32] = S3_d[1152-((36- 8)*32) +: 32] ^ S3_d[1152-((36-30)*32) +: 32];

		S4_d = S3_q;
		S4_d[799:768] = S4[127:96];
		S4_d[831:800] = S4[95:64];
		S4_d[863:832] = S4[63:32];
		S4_d[895:864] = S4[31:0];
		
	end

	always @ (posedge clk) begin

		S0_q <= S0_d;
		S1_q <= S1_d;
		S2_q <= S2_d;
		S3_q <= S3_d;
		S4_q <= S4_d;

	end

endmodule


module close_1 (
	input clk,
	input [1151:0] S,
	output [1151:0] O
);

	wire [127:0] S1;

	reg [1151:0] S0_d, S0_q, S1_d, S1_q;

	smix smix0(S0_q[1152-((36-0)*32) +: 32], S0_q[1152-((36-1)*32) +: 32], S0_q[1152-((36-2)*32) +: 32], S0_q[1152-((36-3)*32) +: 32], S1);
	
	assign O = S1_q;

	always @ (*) begin
	
		S0_d = { S[1055:0], S[1151:1056] };

		// CMIX36
		S0_d[1152-((36-0)*32) +: 32] = S0_d[1152-((36-0)*32) +: 32] ^ S0_d[1152-((36-4)*32) +: 32];
		S0_d[1152-((36-1)*32) +: 32] = S0_d[1152-((36-1)*32) +: 32] ^ S0_d[1152-((36-5)*32) +: 32];
		S0_d[1152-((36-2)*32) +: 32] = S0_d[1152-((36-2)*32) +: 32] ^ S0_d[1152-((36-6)*32) +: 32];
		S0_d[1152-((36-18)*32) +: 32] = S0_d[1152-((36-18)*32) +: 32] ^ S0_d[1152-((36-4)*32) +: 32];
		S0_d[1152-((36-19)*32) +: 32] = S0_d[1152-((36-19)*32) +: 32] ^ S0_d[1152-((36-5)*32) +: 32];
		S0_d[1152-((36-20)*32) +: 32] = S0_d[1152-((36-20)*32) +: 32] ^ S0_d[1152-((36-6)*32) +: 32];

		S1_d = S0_q;
		S1_d[31:0] = S1[127:96];
		S1_d[63:32] = S1[95:64];
		S1_d[95:64] = S1[63:32];
		S1_d[127:96] = S1[31:0];

	end
	
	always @ (posedge clk) begin
	
		S0_q <= S0_d;
		S1_q <= S1_d;

	end

endmodule

module close_2 (
	input clk,
	input [1151:0] S,
	output [1151:0] O
);

	wire [127:0] S1, S2, S3, S4;

	reg [1151:0] S0_d, S1_d, S2_d, S3_d, S4_d;
	reg [1151:0] S0_q, S1_q, S2_q, S3_q, S4_q;
	
	smix smix0 (S0_q[1152-((36-0)*32) +: 32], S0_q[1152-((36-1)*32) +: 32], S0_q[1152-((36-2)*32) +: 32], S0_q[1152-((36-3)*32) +: 32], S1);
	smix smix1 (S1_q[1152-((36-0)*32) +: 32], S1_q[1152-((36-1)*32) +: 32], S1_q[1152-((36-2)*32) +: 32], S1_q[1152-((36-3)*32) +: 32], S2);
	smix smix2 (S2_q[1152-((36-0)*32) +: 32], S2_q[1152-((36-1)*32) +: 32], S2_q[1152-((36-2)*32) +: 32], S2_q[1152-((36-3)*32) +: 32], S3);
	smix smix3 (S3_q[1152-((36-0)*32) +: 32], S3_q[1152-((36-1)*32) +: 32], S3_q[1152-((36-2)*32) +: 32], S3_q[1152-((36-3)*32) +: 32], S4);
	
	assign O = S4_q;
	
	always @ (*) begin
	
		S0_d = S;

		S0_d[1152-((36-4)*32) +: 32] = S0_d[1152-((36-4)*32) +: 32] ^ S0_d[1152-((36-0)*32) +: 32];
		S0_d[1152-((36-9)*32) +: 32] = S0_d[1152-((36-9)*32) +: 32] ^ S0_d[1152-((36-0)*32) +: 32];
		S0_d[1152-((36-18)*32) +: 32] = S0_d[1152-((36-18)*32) +: 32] ^ S0_d[1152-((36-0)*32) +: 32];
		S0_d[1152-((36-27)*32) +: 32] = S0_d[1152-((36-27)*32) +: 32] ^ S0_d[1152-((36-0)*32) +: 32];
		S0_d = { S0_d[863:0], S0_d[1151:864] };

		S1_d = S0_q;
		S1_d[31:0] = S1[127:96];
		S1_d[63:32] = S1[95:64];
		S1_d[95:64] = S1[63:32];
		S1_d[127:96] = S1[31:0];

		S1_d[1152-((36-4)*32) +: 32] = S1_d[1152-((36-4)*32) +: 32] ^ S1_d[1152-((36-0)*32) +: 32];
		S1_d[1152-((36-10)*32) +: 32] = S1_d[1152-((36-10)*32) +: 32] ^ S1_d[1152-((36-0)*32) +: 32];
		S1_d[1152-((36-18)*32) +: 32] = S1_d[1152-((36-18)*32) +: 32] ^ S1_d[1152-((36-0)*32) +: 32];
		S1_d[1152-((36-27)*32) +: 32] = S1_d[1152-((36-27)*32) +: 32] ^ S1_d[1152-((36-0)*32) +: 32];
		S1_d = { S1_d[863:0], S1_d[1151:864] };

		S2_d = S1_q;
		S2_d[31:0] = S2[127:96];
		S2_d[63:32] = S2[95:64];
		S2_d[95:64] = S2[63:32];
		S2_d[127:96] = S2[31:0];

		S2_d[1152-((36-4)*32) +: 32] = S2_d[1152-((36-4)*32) +: 32] ^ S2_d[1152-((36-0)*32) +: 32];
		S2_d[1152-((36-10)*32) +: 32] = S2_d[1152-((36-10)*32) +: 32] ^ S2_d[1152-((36-0)*32) +: 32];
		S2_d[1152-((36-19)*32) +: 32] = S2_d[1152-((36-19)*32) +: 32] ^ S2_d[1152-((36-0)*32) +: 32];
		S2_d[1152-((36-27)*32) +: 32] = S2_d[1152-((36-27)*32) +: 32] ^ S2_d[1152-((36-0)*32) +: 32];
		S2_d = { S2_d[863:0], S2_d[1151:864] };

		S3_d = S2_q;
		S3_d[31:0] = S3[127:96];
		S3_d[63:32] = S3[95:64];
		S3_d[95:64] = S3[63:32];
		S3_d[127:96] = S3[31:0];

		S3_d[1152-((36-4)*32) +: 32] = S3_d[1152-((36-4)*32) +: 32] ^ S3_d[1152-((36-0)*32) +: 32];
		S3_d[1152-((36-10)*32) +: 32] = S3_d[1152-((36-10)*32) +: 32] ^ S3_d[1152-((36-0)*32) +: 32];
		S3_d[1152-((36-19)*32) +: 32] = S3_d[1152-((36-19)*32) +: 32] ^ S3_d[1152-((36-0)*32) +: 32];
		S3_d[1152-((36-28)*32) +: 32] = S3_d[1152-((36-28)*32) +: 32] ^ S3_d[1152-((36-0)*32) +: 32];
		S3_d = { S3_d[895:0], S3_d[1151:896] };

		S4_d = S3_q;
		S4_d[31:0] = S4[127:96];
		S4_d[63:32] = S4[95:64];
		S4_d[95:64] = S4[63:32];
		S4_d[127:96] = S4[31:0];

	end

	always @ (posedge clk) begin

		S0_q <= S0_d;
		S1_q <= S1_d;
		S2_q <= S2_d;
		S3_q <= S3_d;
		S4_q <= S4_d;

	end

endmodule

